 library IEEE;
 use IEEE.STD_LOGIC_1164.all;
 use IEEE.NUMERIC_STD.ALL;

 package mat_pak is
	  type matrix  is array (natural range <>, natural range <>) of std_logic;                    
 end mat_pak;
